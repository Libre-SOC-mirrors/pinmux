/* ==== define the AXI Addresses ==== */
{0}


