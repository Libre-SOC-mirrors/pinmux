`define ADDR 32
`define DATA 64
`define USERSPACE 0
