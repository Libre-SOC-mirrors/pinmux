`define ADDR 32
`define DATA 64
`define USERSPACE 0
`define PADDR 32
`define Reg_width 32
