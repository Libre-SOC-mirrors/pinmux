/*====== Fast peripherals Memory Map ======= */
{0}
